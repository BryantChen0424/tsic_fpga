/*
 *  icebreaker examples - Async uart mirror using pll
 *
 *  Copyright (C) 2018 Piotr Esden-Tempski <piotr@esden.net>
 *
 *  Modified work
 *  Copyright (C) 2025 Bryant Chen <bryant90424@gmail.com>
 *
 *  Permission to use, copy, modify, and/or distribute this software for any
 *  purpose with or without fee is hereby granted, provided that the above
 *  copyright notice and this permission notice appear in all copies.
 *
 *  THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
 *  WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
 *  MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
 *  ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
 *  WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
 *  ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
 *  OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 *
 */

module top (
	input  clk,
	input RX,
    output reg TX
);

function integer log2(input integer v); begin
	log2 = 0;
	while(v >> log2) log2 = log2 + 1;
end endfunction

localparam WIDTH = 8;
localparam LEN = 256;

localparam TXSTR_BASE = LEN/2;

reg [log2(LEN-1):0] addr;
reg [WIDTH-1:0] din;
wire [WIDTH-1:0] dout;
reg we;

bram #(WIDTH, LEN) mem (
    .clk(clk),
    .addr(addr),
    .din(din),
    .dout(dout),
    .we(we)
);

wire rx_ready;
wire [7:0] rx_data;

uart_rx #(12_000_000, 115200) urx (
    .clk(clk),
    .rx(RX),
    .rx_ready(rx_ready),
    .rx_data(rx_data)
);

reg tx_start;
reg [7:0] tx_data;
wire tx_busy;

uart_tx #(12_000_000, 115200) utx (
    .clk(clk),
    .tx_start(tx_start),
    .tx_data(tx_data),
    .tx(TX),
    .tx_busy(tx_busy)
);

reg echo_rx_ready;
reg [7:0] echo_rx_data;

wire echo_tx_start;
wire [7:0] echo_tx_data;
reg echo_tx_busy;

reg echo_get_a_cmd = 0;
wire echo_idle;

uart_echo_unit #(12_000_000, 115200) ueu (
    .clk(clk),

    .rx_data(echo_rx_data),
    .rx_ready(echo_rx_ready),

    .tx_start(echo_tx_start),
    .tx_data(echo_tx_data),
    .tx_busy(echo_tx_busy),

    .get_a_cmd(echo_get_a_cmd),
    .idle(echo_idle)
);

////////////////

localparam S_rst = 0;
localparam S_Rp  = 1;
localparam S_R   = 2;
localparam S_Rf  = 3;
localparam S_NL  = 4;
localparam S_T   = 5;

reg [3:0] S = S_rst;

reg [log2(LEN-1):0] rx_line_len = 0;
reg [log2(LEN-1):0] tx_line_len = 0;

reg resp_tx_start = 0;
reg [7:0] resp_tx_data = 0;
reg resp_tx_busy;

reg nl2tx_flag = 0;
reg tx_flag = 0;

////////////////

always @(*) begin
    echo_tx_busy = tx_busy;
    resp_tx_busy = tx_busy;

    echo_rx_data = rx_data;
    echo_rx_ready = rx_ready;
    case (S)
        S_Rp: begin
            tx_start = 0;
            tx_data = 0;
        end
        S_R: begin
            tx_start = echo_tx_start;
            tx_data = echo_tx_data;
        end
        S_Rf: begin
            tx_start = echo_tx_start;
            tx_data = echo_tx_data;
        end
        S_NL: begin
            tx_start = 0;
            tx_data = 0;
        end
        S_T: begin
            tx_start = resp_tx_start;
            tx_data = resp_tx_data;
        end
        default: begin
            tx_start = 0;
            tx_data = 0;
        end
    endcase
end

////////////////

reg [15:0] rst_cnt;

always @(posedge clk) begin
    rst_cnt <= rst_cnt + 1;
    case (S)
        S_rst: begin
            if (rst_cnt[15]) begin
                S <= S_Rp;
            end
        end
        S_Rp: begin
            echo_get_a_cmd <= 1; 
            S <= S_R;
        end
        S_R: begin
            echo_get_a_cmd <= 0;
            if (rx_ready) begin
                addr <= rx_line_len;
                din <= echo_rx_data;
                we <= 1;

                rx_line_len <= rx_line_len + 1;
            end
            else begin
                din <= 0;
                we <= 0;
            end

            if (din == "\r" || din == "\n") begin
                S <= S_Rf;
            end

            tx_line_len <= 0;
        end
        S_Rf: begin
            if (echo_idle) begin
                S <= S_NL;
            end
        end
        S_NL: begin
            if (tx_line_len == 30) begin
                addr <= TXSTR_BASE;
                din <= 0;
                we <= 0;

                nl2tx_flag <= 0;
                S <= S_T;
            end
            else if (tx_line_len == 29) begin
                addr <= tx_line_len + TXSTR_BASE;
                din <= "\r";
                we <= 1;

                tx_line_len <= tx_line_len + 1;
            end
            else if (tx_line_len == 28) begin
                addr <= tx_line_len + TXSTR_BASE;
                din <= "\n";
                we <= 1;

                tx_line_len <= tx_line_len + 1;
            end
            else begin
                addr <= tx_line_len + TXSTR_BASE;
                din <= tx_line_len + 64;
                we <= 1;

                tx_line_len <= tx_line_len + 1;
            end
        end
        S_T: begin
            if (~nl2tx_flag) begin
                nl2tx_flag <= 1;
            end
            else begin
                if (~tx_flag) begin
                    resp_tx_start <= 1;
                    resp_tx_data <= dout;
                    tx_flag <= 1;

                    addr <= addr + 1;
                end
                else begin
                    if (resp_tx_start) begin
                        resp_tx_start <= 0;
                        resp_tx_data <= 0;
                    end
                    else if (~resp_tx_busy) begin
                        tx_flag <= 0;
                        if (addr == tx_line_len + TXSTR_BASE) begin
                            S <= S_Rp;
                        end
                    end
                end
            end
        end
        default: begin
            
        end
    endcase
    
end

endmodule
