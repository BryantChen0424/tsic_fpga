module top (
    input  wire clk,

    input RX,
    output TX,

    output wire oled_cs,
    output wire oled_clk,
    output wire oled_mosi,
    output wire oled_dc,
    output wire reset
);

localparam X_MAX = 160;
localparam Y_MAX = 80;

localparam CLK_FREQ = 12000000;
localparam BAUD = 115200;

function integer log2(input integer v); begin
	log2 = 0;
	while(v >> log2) log2 = log2 + 1;
end endfunction

wire rx_ready;
wire [7:0] rx_data;

uart_rx #(CLK_FREQ, BAUD) urx (
    .clk(clk),
    .rx(RX),
    .rx_ready(rx_ready),
    .rx_data(rx_data)
);

reg tx_start;
reg [7:0] tx_data;
wire tx_busy;

uart_tx #(CLK_FREQ, BAUD) utx (
    .clk(clk),
    .tx_start(tx_start),
    .tx_data(tx_data),
    .tx(TX),
    .tx_busy(tx_busy)
);

uart_echo_unit #(CLK_FREQ, BAUD) ueu (
    .clk(clk),

    .rx_data(rx_data),
    .rx_ready(rx_ready),

    .tx_start(tx_start),
    .tx_data(tx_data),
    .tx_busy(tx_busy),

    .en(1),
    .idle()
);

reg [15:0] color;
wire [7:0] x;
wire [6:0] y;
wire next_pixel;

st7735  driver (
    .clk(clk),
    .x(x),
    .y(y),
    .color(color),
    .next_pixel(next_pixel),

    .oled_cs(oled_cs),
    .oled_clk(oled_clk),
    .oled_mosi(oled_mosi),
    .oled_dc(oled_dc),
    .reset(reset)
);

localparam SRC_BASE = X_MAX * Y_MAX;
localparam WIDTH = 4;
localparam LEN = SRC_BASE + 2000;

reg [log2(LEN-1):0] addr;
reg [WIDTH-1:0] din;
wire [WIDTH-1:0] dout;
reg we;

bram #(WIDTH, LEN) mem (
    .clk(clk),
    .addr(addr),
    .din(din),
    .dout(dout),
    .we(we)
);

localparam RND_WIDTH = 8;

reg rndg_en = 1;
reg rndg_load_seed = 1;
reg [RND_WIDTH-1:0] rndg_seed = 0;
wire [RND_WIDTH-1:0] rndg_rnd;

rnd_gen #(RND_WIDTH) rndg (
    .clk(clk),
    .rst_n(reset),
    .en(rndg_en),        
    .load_seed(rndg_load_seed), 
    .seed(rndg_seed),      
    .rnd(rndg_rnd)        
);

reg [15:0] digits_sel = 0;

localparam S_UPDATE = 0;
localparam S_DISPLAY = 1;

reg S = S_DISPLAY;

reg u_update;
wire u_done;

wire [log2(LEN-1):0] u_addr;
wire [WIDTH-1:0] u_din;
reg [WIDTH-1:0] u_dout;
wire u_we;

display_buf_updater #(LEN, WIDTH, X_MAX, Y_MAX) dbu (
    .clk(clk),
    .rst_n(reset),

    .update(u_update),
    .done(u_done),

    .addr(u_addr),
    .din(u_din),
    .dout(u_dout),
    .we(u_we),

    .digits_sel(digits_sel)
);

always @(*) begin
    u_dout = dout;
    case (S)
        S_UPDATE: begin
            addr = u_addr;
            din = u_din;
            we = u_we;
        end 
        S_DISPLAY: begin
            addr = y * 160 + x;
            din = 0;
            we = 0;
        end
    endcase
end

always @(posedge clk) begin
    if (~reset) begin
        digits_sel <= 0;
        seed_flag <= 0;

        S <= S_DISPLAY;
    end
    else begin
        case (S)
            S_UPDATE: begin
                u_update <= 0;
                if (u_done) begin
                    S <= S_DISPLAY;
                end
            end
            S_DISPLAY: begin
                if (next_pixel) begin
                    color <= {
                        {dout, 1'b0},
                        {dout, 2'b0},
                        {dout, 1'b0}
                    };
                end
                if (rx_ready && ~seed_flag) begin
                    digits_sel <= (rndg_seed * 10) >> 8;
                    rndg_load_seed <= 1;
                    u_update <= 1;
                    S <= S_UPDATE;
                end
                else if (rx_ready && seed_flag) begin
                    digits_sel <= (rndg_rnd * 10) >> 8;
                    u_update <= 1;
                    S <= S_UPDATE;
                end
                else begin
                    rndg_load_seed <= 0;
                end
            end
        endcase

        rndg_seed <= rndg_seed + 1;
        seed_flag <= seed_flag | rx_ready;
    end
end

endmodule

